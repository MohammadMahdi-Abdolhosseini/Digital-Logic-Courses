`timescale 1ns/1ns
module barrelShifter16Bit (input [15:0] A, input [3:0] S, output [15:0] SHO);
	
	wire [15:0] J1,J2,J3,J4,J5,J6,J7,J8,J9,J10,J11,J12,J13,J14,J15,J16;
	assign J1 = {A[14],  A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15]};
	assign J2 = {A[13],  A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14]};
	assign J3 = {A[12],  A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13]};
	assign J4 = {A[11],  A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12]};
	assign J5 = {A[10],  A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11]};
	assign J6 = {A[9],   A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10]};
	assign J7 = {A[8],   A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9]};
	assign J8 = {A[7],   A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8]};
	assign J9 = {A[6],   A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7]};
	assign J10 = {A[5],  A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6]};
	assign J11 = {A[4],  A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5]};
	assign J12 = {A[3],  A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4]};
	assign J13 = {A[2],  A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3]};
	assign J14 = {A[1],  A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2]};
	assign J15 = {A[0],  A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1]};
	assign J16 = {A[15], A[14], A[13], A[12], A[11], A[10], A[9],  A[8],  A[7],  A[6],  A[5],  A[4],  A[3],  A[2],  A[1],  A[0]};
	mux16to1 M1(J1, S, SHO[15]);
	mux16to1 M2(J2, S, SHO[14]);
	mux16to1 M3(J3, S, SHO[13]);
	mux16to1 M4(J4, S, SHO[12]);
	mux16to1 M5(J5, S, SHO[11]);
	mux16to1 M6(J6, S, SHO[10]);
	mux16to1 M7(J7, S, SHO[9]);
	mux16to1 M8(J8, S, SHO[8]);
	mux16to1 M9(J9, S, SHO[7]);
	mux16to1 M10(J10, S, SHO[6]);
	mux16to1 M11(J11, S, SHO[5]);
	mux16to1 M12(J12, S, SHO[4]);
	mux16to1 M13(J13, S, SHO[3]);
	mux16to1 M14(J14, S, SHO[2]);
	mux16to1 M15(J15, S, SHO[1]);
	mux16to1 M16(J16, S, SHO[0]);
	
endmodule

